module NotGate(
    input  a,
    output y
);
    assign y = ~a;
endmodule